magic
tech scmos
timestamp 1580705360
<< nwell >>
rect -8 46 86 66
<< polysilicon >>
rect 8 62 10 65
rect 38 62 40 65
rect 68 62 70 65
rect 8 8 10 50
rect 38 8 40 50
rect 68 8 70 50
rect 8 -7 10 -4
rect 38 -7 40 -4
rect 68 -7 70 -4
<< ndiffusion >>
rect -4 4 8 8
rect -4 0 0 4
rect 4 0 8 4
rect -4 -4 8 0
rect 10 4 22 8
rect 10 0 14 4
rect 18 0 22 4
rect 10 -4 22 0
rect 26 4 38 8
rect 26 0 30 4
rect 34 0 38 4
rect 26 -4 38 0
rect 40 4 52 8
rect 40 0 44 4
rect 48 0 52 4
rect 40 -4 52 0
rect 56 4 68 8
rect 56 0 60 4
rect 64 0 68 4
rect 56 -4 68 0
rect 70 4 82 8
rect 70 0 74 4
rect 78 0 82 4
rect 70 -4 82 0
<< pdiffusion >>
rect -4 58 8 62
rect -4 54 0 58
rect 4 54 8 58
rect -4 50 8 54
rect 10 50 38 62
rect 40 50 68 62
rect 70 58 82 62
rect 70 54 74 58
rect 78 54 82 58
rect 70 50 82 54
<< metal1 >>
rect 0 78 78 82
rect 0 74 4 78
rect 8 74 34 78
rect 38 74 64 78
rect 68 74 78 78
rect 0 70 78 74
rect 0 58 4 70
rect 0 50 4 54
rect 74 58 78 62
rect 74 32 78 54
rect 0 28 4 32
rect 30 28 34 32
rect 60 28 64 32
rect 74 28 86 32
rect 74 20 78 28
rect 14 16 78 20
rect 0 4 4 8
rect 0 -11 4 0
rect 14 4 18 16
rect 14 -4 18 0
rect 30 4 34 8
rect 30 -11 34 0
rect 44 4 48 16
rect 44 -4 48 0
rect 60 4 64 8
rect 60 -11 64 0
rect 74 4 78 16
rect 74 -4 78 0
rect 0 -15 78 -11
rect 0 -19 4 -15
rect 8 -19 34 -15
rect 38 -19 64 -15
rect 68 -19 78 -15
rect 0 -23 78 -19
<< ntransistor >>
rect 8 -4 10 8
rect 38 -4 40 8
rect 68 -4 70 8
<< ptransistor >>
rect 8 50 10 62
rect 38 50 40 62
rect 68 50 70 62
<< polycontact >>
rect 4 28 8 32
rect 34 28 38 32
rect 64 28 68 32
<< ndcontact >>
rect 0 0 4 4
rect 14 0 18 4
rect 30 0 34 4
rect 44 0 48 4
rect 60 0 64 4
rect 74 0 78 4
<< pdcontact >>
rect 0 54 4 58
rect 74 54 78 58
<< psubstratepcontact >>
rect 4 74 8 78
rect 34 74 38 78
rect 64 74 68 78
<< nsubstratencontact >>
rect 4 -19 8 -15
rect 34 -19 38 -15
rect 64 -19 68 -15
<< labels >>
rlabel metal1 0 70 78 82 1 vdd
rlabel metal1 0 -23 78 -11 1 gnd
rlabel metal1 0 28 8 32 1 a
rlabel metal1 30 28 38 32 1 b
rlabel metal1 60 28 68 32 1 c
rlabel metal1 78 28 86 32 7 out
<< end >>
