magic
tech scmos
timestamp 1580703964
<< nwell >>
rect -8 36 40 56
<< polysilicon >>
rect 8 52 10 55
rect 22 52 24 55
rect 8 8 10 40
rect 22 8 24 40
rect 8 -7 10 -4
rect 22 -7 24 -4
<< ndiffusion >>
rect -4 4 8 8
rect -4 0 0 4
rect 4 0 8 4
rect -4 -4 8 0
rect 10 4 22 8
rect 10 0 14 4
rect 18 0 22 4
rect 10 -4 22 0
rect 24 4 36 8
rect 24 0 28 4
rect 32 0 36 4
rect 24 -4 36 0
<< pdiffusion >>
rect -4 48 8 52
rect -4 44 0 48
rect 4 44 8 48
rect -4 40 8 44
rect 10 40 22 52
rect 24 48 36 52
rect 24 44 28 48
rect 32 44 36 48
rect 24 40 36 44
<< metal1 >>
rect 0 71 32 75
rect 0 67 4 71
rect 8 67 14 71
rect 18 67 24 71
rect 28 67 32 71
rect 0 63 32 67
rect 0 48 4 63
rect 0 40 4 44
rect 28 48 32 52
rect 0 27 4 31
rect 28 25 32 44
rect 14 21 40 25
rect 0 4 4 8
rect 0 -11 4 0
rect 14 4 18 21
rect 28 13 32 17
rect 14 -4 18 0
rect 28 4 32 8
rect 28 -11 32 0
rect 0 -15 32 -11
rect 0 -19 4 -15
rect 8 -19 14 -15
rect 18 -19 24 -15
rect 28 -19 32 -15
rect 0 -23 32 -19
<< ntransistor >>
rect 8 -4 10 8
rect 22 -4 24 8
<< ptransistor >>
rect 8 40 10 52
rect 22 40 24 52
<< polycontact >>
rect 4 27 8 31
rect 24 13 28 17
<< ndcontact >>
rect 0 0 4 4
rect 14 0 18 4
rect 28 0 32 4
<< pdcontact >>
rect 0 44 4 48
rect 28 44 32 48
<< psubstratepcontact >>
rect 4 67 8 71
rect 14 67 18 71
rect 24 67 28 71
<< nsubstratencontact >>
rect 4 -19 8 -15
rect 14 -19 18 -15
rect 24 -19 28 -15
<< labels >>
rlabel metal1 0 63 32 75 1 vdd
rlabel metal1 0 -23 32 -11 1 gnd
rlabel metal1 24 13 32 17 1 b
rlabel metal1 0 27 8 31 1 a
rlabel metal1 32 21 40 25 7 out
<< end >>
