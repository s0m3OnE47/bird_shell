magic
tech scmos
timestamp 1581044992
<< nwell >>
rect -8 -8 86 12
<< polysilicon >>
rect 8 8 10 11
rect 38 8 40 11
rect 68 8 70 12
rect 8 -28 10 -4
rect 38 -28 40 -4
rect 68 -28 70 -4
rect 8 -43 10 -40
rect 38 -43 40 -40
rect 68 -42 70 -40
<< ndiffusion >>
rect -4 -32 8 -28
rect -4 -36 0 -32
rect 4 -36 8 -32
rect -4 -40 8 -36
rect 10 -40 38 -28
rect 40 -40 68 -28
rect 70 -32 82 -28
rect 70 -36 74 -32
rect 78 -36 82 -32
rect 70 -40 82 -36
<< pdiffusion >>
rect -4 4 8 8
rect -4 0 0 4
rect 4 0 8 4
rect -4 -4 8 0
rect 10 4 22 8
rect 10 0 14 4
rect 18 0 22 4
rect 10 -4 22 0
rect 26 4 38 8
rect 26 0 30 4
rect 34 0 38 4
rect 26 -4 38 0
rect 40 4 52 8
rect 40 0 44 4
rect 48 0 52 4
rect 40 -4 52 0
rect 56 4 68 8
rect 56 0 60 4
rect 64 0 68 4
rect 56 -4 68 0
rect 70 4 82 8
rect 70 0 74 4
rect 78 0 82 4
rect 70 -4 82 0
<< metal1 >>
rect 0 24 64 28
rect 0 20 4 24
rect 8 20 26 24
rect 30 20 56 24
rect 60 20 64 24
rect 0 16 64 20
rect 0 4 4 16
rect 0 -4 4 0
rect 14 4 18 8
rect 14 -14 18 0
rect 30 4 34 16
rect 30 -4 34 0
rect 44 4 48 8
rect 44 -14 48 0
rect 60 4 64 16
rect 60 -4 64 0
rect 74 4 78 8
rect 74 -14 78 0
rect 14 -18 86 -14
rect 0 -25 4 -21
rect 30 -25 34 -21
rect 60 -25 64 -21
rect 0 -32 4 -28
rect 0 -48 4 -36
rect 74 -32 78 -18
rect 74 -40 78 -36
rect 0 -52 64 -48
rect 0 -56 4 -52
rect 8 -56 26 -52
rect 30 -56 56 -52
rect 60 -56 64 -52
rect 0 -60 64 -56
<< ntransistor >>
rect 8 -40 10 -28
rect 38 -40 40 -28
rect 68 -40 70 -28
<< ptransistor >>
rect 8 -4 10 8
rect 38 -4 40 8
rect 68 -4 70 8
<< polycontact >>
rect 4 -25 8 -21
rect 34 -25 38 -21
rect 64 -25 68 -21
<< ndcontact >>
rect 0 -36 4 -32
rect 74 -36 78 -32
<< pdcontact >>
rect 0 0 4 4
rect 14 0 18 4
rect 30 0 34 4
rect 44 0 48 4
rect 60 0 64 4
rect 74 0 78 4
<< psubstratepcontact >>
rect 4 20 8 24
rect 26 20 30 24
rect 56 20 60 24
<< nsubstratencontact >>
rect 4 -56 8 -52
rect 26 -56 30 -52
rect 56 -56 60 -52
<< labels >>
rlabel metal1 0 -60 64 -48 1 gnd
rlabel metal1 0 16 64 28 1 vcc
rlabel metal1 0 -25 8 -21 1 a
rlabel metal1 30 -25 38 -21 1 b
rlabel metal1 60 -25 68 -21 1 c
rlabel metal1 78 -18 86 -14 7 out
<< end >>
