magic
tech scmos
timestamp 1581047204
<< nwell >>
rect -8 -8 54 12
<< polysilicon >>
rect 8 8 10 11
rect 22 8 24 11
rect 36 8 38 11
rect 8 -32 10 -4
rect 22 -32 24 -4
rect 36 -32 38 -4
rect 8 -47 10 -44
rect 22 -47 24 -44
rect 36 -47 38 -44
<< ndiffusion >>
rect -4 -36 8 -32
rect -4 -40 0 -36
rect 4 -40 8 -36
rect -4 -44 8 -40
rect 10 -44 22 -32
rect 24 -44 36 -32
rect 38 -36 50 -32
rect 38 -40 42 -36
rect 46 -40 50 -36
rect 38 -44 50 -40
<< pdiffusion >>
rect -4 4 8 8
rect -4 0 0 4
rect 4 0 8 4
rect -4 -4 8 0
rect 10 4 22 8
rect 10 0 14 4
rect 18 0 22 4
rect 10 -4 22 0
rect 24 4 36 8
rect 24 0 28 4
rect 32 0 36 4
rect 24 -4 36 0
rect 38 4 50 8
rect 38 0 42 4
rect 46 0 50 4
rect 38 -4 50 0
<< metal1 >>
rect 0 24 40 28
rect 0 20 4 24
rect 8 20 18 24
rect 22 20 32 24
rect 36 20 40 24
rect 0 16 40 20
rect 0 4 4 16
rect 0 -4 4 0
rect 14 4 18 8
rect 42 4 46 8
rect 14 -15 18 0
rect 42 -15 46 0
rect 14 -19 46 -15
rect 42 -23 46 -19
rect 0 -27 4 -23
rect 14 -27 18 -23
rect 28 -27 32 -23
rect 42 -27 54 -23
rect 0 -36 4 -32
rect 0 -51 4 -40
rect 42 -36 46 -27
rect 42 -44 46 -40
rect 0 -55 40 -51
rect 0 -59 4 -55
rect 8 -59 18 -55
rect 22 -59 32 -55
rect 36 -59 40 -55
rect 0 -63 40 -59
<< ntransistor >>
rect 8 -44 10 -32
rect 22 -44 24 -32
rect 36 -44 38 -32
<< ptransistor >>
rect 8 -4 10 8
rect 22 -4 24 8
rect 36 -4 38 8
<< polycontact >>
rect 4 -27 8 -23
rect 18 -27 22 -23
rect 32 -27 36 -23
<< ndcontact >>
rect 0 -40 4 -36
rect 42 -40 46 -36
<< pdcontact >>
rect 0 0 4 4
rect 14 0 18 4
rect 28 0 32 4
rect 42 0 46 4
<< psubstratepcontact >>
rect 4 20 8 24
rect 18 20 22 24
rect 32 20 36 24
<< nsubstratencontact >>
rect 4 -59 8 -55
rect 18 -59 22 -55
rect 32 -59 36 -55
<< labels >>
rlabel metal1 0 16 40 28 1 vdd
rlabel metal1 0 -63 40 -51 1 gnd
rlabel metal1 0 -27 8 -23 1 a
rlabel metal1 14 -27 22 -23 1 v
rlabel metal1 28 -27 36 -23 1 b
rlabel metal1 46 -27 54 -23 7 out
<< end >>
